localparam BP_TWOBIT       = (32'd0);
localparam BP_GSHARE       = (32'd1);
localparam BP_GLOBAL       = (32'd2);
localparam BP_GSHARE_BASIC = (32'd3);
localparam BP_GLOBAL_BASIC = (32'd4);
localparam BP_LOCAL_BASIC  = (32'd5);
localparam BP_LOCAL_AHEAD  = (32'd6);
localparam BP_LOCAL_REPAIR = (32'd7);
